*** SPICE deck for cell xor_sim{lay} from library project_1
*** Created on Thu Oct 24, 2024 14:30:56
*** Last revised on Thu Oct 24, 2024 14:34:11
*** Written on Thu Oct 24, 2024 14:34:27 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project_1__xor FROM CELL xor{lay}
.SUBCKT project_1__xor A B gnd out vdd
Mnmos@7 net@7 net@70 gnd gnd NMOS L=0.35U W=1.75U AS=9.188P AD=1.302P PS=19.775U PD=3.238U
Mnmos@11 out net@94 net@7 gnd NMOS L=0.35U W=1.75U AS=1.302P AD=1.493P PS=3.238U PD=3.456U
Mnmos@12 gnd A net@11 gnd NMOS L=0.35U W=1.75U AS=1.608P AD=9.188P PS=3.588U PD=19.775U
Mnmos@13 net@11 B out gnd NMOS L=0.35U W=1.75U AS=1.493P AD=1.608P PS=3.456U PD=3.588U
Mnmos@14 net@70 B gnd gnd NMOS L=0.35U W=1.75U AS=9.188P AD=2.45P PS=19.775U PD=6.3U
Mnmos@15 gnd A net@94 gnd NMOS L=0.35U W=1.75U AS=1.991P AD=9.188P PS=5.775U PD=19.775U
Mpmos@7 out net@70 net@0 vdd PMOS L=0.35U W=1.75U AS=1.991P AD=1.493P PS=4.9U PD=3.456U
Mpmos@9 net@0 net@94 out vdd PMOS L=0.35U W=1.75U AS=1.493P AD=1.991P PS=3.456U PD=4.9U
Mpmos@10 net@0 A vdd vdd PMOS L=0.35U W=1.75U AS=8.843P AD=1.991P PS=18.506U PD=4.9U
Mpmos@11 vdd B net@0 vdd PMOS L=0.35U W=1.75U AS=1.991P AD=8.843P PS=4.9U PD=18.506U
Mpmos@12 net@70 B vdd vdd PMOS L=0.35U W=1.75U AS=8.843P AD=2.45P PS=18.506U PD=6.3U
Mpmos@13 vdd A net@94 vdd PMOS L=0.35U W=1.75U AS=1.991P AD=8.843P PS=5.775U PD=18.506U
.ENDS project_1__xor

*** TOP LEVEL CELL: xor_sim{lay}
Xxor@0 A B gnd out vdd project_1__xor

* Spice Code nodes in cell cell 'xor_sim{lay}'
vdd vdd 0 dc 5 
va A 0 pulse 0 5 0 2n 3n 250n 500n 
vb B 0 pulse 0 5 0 2n 3n 125n 250n 
cload out 0 250fF
.tran 0 1u 
.include D:\C5_models.txt
.END

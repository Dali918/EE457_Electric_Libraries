*** SPICE deck for cell xor{sch} from library project_1
*** Created on Wed Oct 16, 2024 20:40:51
*** Last revised on Sat Oct 19, 2024 18:49:33
*** Written on Sat Oct 19, 2024 18:49:39 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project_1__inv_10_10 FROM CELL inv_10_10{sch}
.SUBCKT project_1__inv_10_10 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 out in vdd vdd PMOS L=0.35U W=1.75U
.ENDS project_1__inv_10_10

.global gnd vdd

*** TOP LEVEL CELL: xor{sch}
Mnmos@6 net@194 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@9 net@195 net@224 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@10 net@135 B net@194 gnd NMOS L=0.35U W=1.75U
Mnmos@11 net@135 net@231 net@195 gnd NMOS L=0.35U W=1.75U
Mpmos@9 net@186 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@10 net@135 B net@186 vdd PMOS L=0.35U W=1.75U
Mpmos@11 net@186 net@224 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@12 net@135 net@231 net@186 vdd PMOS L=0.35U W=1.75U
Xinv_10_1@0 net@135 out project_1__inv_10_10
Xinv_20_1@0 A net@231 project_1__inv_10_10
Xinv_20_1@1 B net@224 project_1__inv_10_10
.END

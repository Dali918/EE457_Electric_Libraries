*** SPICE deck for cell 8bit_ripple{sch} from library project_1
*** Created on Sun Oct 20, 2024 23:17:08
*** Last revised on Tue Oct 22, 2024 02:57:58
*** Written on Tue Oct 22, 2024 10:56:05 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project_1__full_adder FROM CELL full_adder{sch}
.SUBCKT project_1__full_adder A B Cin Cout Sout
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@17 Cin net@31 gnd NMOS L=0.35U W=1.75U
Mnmos@1 net@31 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@2 net@31 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@3 net@17 A net@30 gnd NMOS L=0.35U W=1.75U
Mnmos@4 net@30 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@5 net@108 net@17 net@125 gnd NMOS L=0.35U W=1.75U
Mnmos@6 net@125 Cin gnd gnd NMOS L=0.35U W=1.75U
Mnmos@7 net@125 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@8 net@125 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@9 net@108 A net@264 gnd NMOS L=0.35U W=1.75U
Mnmos@10 net@264 B net@263 gnd NMOS L=0.35U W=1.75U
Mnmos@11 net@263 Cin gnd gnd NMOS L=0.35U W=1.75U
Mnmos@12 Cout net@17 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@13 Sout net@108 gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 net@6 Cin vdd vdd PMOS L=0.35U W=1.75U
Mpmos@1 net@83 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@2 net@6 B net@83 vdd PMOS L=0.35U W=1.75U
Mpmos@3 net@17 B net@6 vdd PMOS L=0.35U W=1.75U
Mpmos@4 net@17 A net@6 vdd PMOS L=0.35U W=1.75U
Mpmos@5 net@98 net@17 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@9 net@108 B net@98 vdd PMOS L=0.35U W=1.75U
Mpmos@10 net@108 Cin net@98 vdd PMOS L=0.35U W=1.75U
Mpmos@11 net@108 A net@98 vdd PMOS L=0.35U W=1.75U
Mpmos@12 net@205 B vdd vdd PMOS L=0.35U W=1.75U
Mpmos@13 net@207 Cin net@205 vdd PMOS L=0.35U W=1.75U
Mpmos@14 net@98 A net@207 vdd PMOS L=0.35U W=1.75U
Mpmos@15 Cout net@17 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@16 Sout net@108 vdd vdd PMOS L=0.35U W=1.75U
.ENDS project_1__full_adder

*** SUBCIRCUIT project_1__inv_10_10 FROM CELL inv_10_10{sch}
.SUBCKT project_1__inv_10_10 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 out in vdd vdd PMOS L=0.35U W=1.75U
.ENDS project_1__inv_10_10

*** SUBCIRCUIT project_1__xor FROM CELL xor{sch}
.SUBCKT project_1__xor A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@6 net@194 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@9 net@195 net@292 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@10 out B net@194 gnd NMOS L=0.35U W=1.75U
Mnmos@11 out net@289 net@195 gnd NMOS L=0.35U W=1.75U
Mpmos@9 net@186 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@10 out net@289 net@186 vdd PMOS L=0.35U W=1.75U
Mpmos@11 net@186 B vdd vdd PMOS L=0.35U W=1.75U
Mpmos@12 out net@292 net@186 vdd PMOS L=0.35U W=1.75U
Xinv_20_1@0 B net@292 project_1__inv_10_10
Xinv_20_1@1 A net@289 project_1__inv_10_10
.ENDS project_1__xor

.global gnd vdd

*** TOP LEVEL CELL: 8bit_ripple{sch}
Xfull_adder_[0] A[0] Bx[0] Cin carry[0] Sout[0] project_1__full_adder
Xfull_adder_[1] A[1] Bx[1] carry[0] carry[1] Sout[1] project_1__full_adder
Xfull_adder_[2] A[2] Bx[2] carry[1] carry[2] Sout[2] project_1__full_adder
Xfull_adder_[3] A[3] Bx[3] carry[2] carry[3] Sout[3] project_1__full_adder
Xfull_adder_[4] A[4] Bx[4] carry[3] carry[4] Sout[4] project_1__full_adder
Xfull_adder_[5] A[5] Bx[5] carry[4] carry[5] Sout[5] project_1__full_adder
Xfull_adder_[6] A[6] Bx[6] carry[5] carry[6] Sout[6] project_1__full_adder
Xfull_adder_[7] A[7] Bx[7] carry[6] Cout Sout[7] project_1__full_adder
Xxor[0] B[0] Cin Bx[0] project_1__xor
Xxor[1] B[1] Cin Bx[1] project_1__xor
Xxor[2] B[2] Cin Bx[2] project_1__xor
Xxor[3] B[3] Cin Bx[3] project_1__xor
Xxor[4] B[4] Cin Bx[4] project_1__xor
Xxor[5] B[5] Cin Bx[5] project_1__xor
Xxor[6] B[6] Cin Bx[6] project_1__xor
Xxor[7] B[7] Cin Bx[7] project_1__xor
.END

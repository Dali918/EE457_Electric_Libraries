*** SPICE deck for cell NAND_sim{lay} from library tutorial_4
*** Created on Tue Oct 15, 2024 23:59:47
*** Last revised on Wed Oct 16, 2024 00:14:52
*** Written on Wed Oct 16, 2024 00:19:38 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT tutorial_4__NAND_2 FROM CELL NAND_2{lay}
.SUBCKT tutorial_4__NAND_2 A AnandB B gnd vdd
Mnmos@1 net@35 B gnd gnd NMOS L=0.35U W=1.75U AS=6.584P AD=0.689P PS=18.025U PD=2.537U
Mnmos@2 AnandB A net@35 gnd NMOS L=0.35U W=1.75U AS=0.689P AD=1.48P PS=2.537U PD=4.025U
Mpmos@1 vdd B AnandB vdd PMOS L=0.35U W=1.75U AS=1.48P AD=4.211P PS=4.025U PD=11.813U
Mpmos@2 AnandB A vdd vdd PMOS L=0.35U W=1.75U AS=4.211P AD=1.48P PS=11.813U PD=4.025U
.ENDS tutorial_4__NAND_2

*** TOP LEVEL CELL: NAND_sim{lay}
XNAND_2@1 in out vdd gnd vdd tutorial_4__NAND_2

* Spice Code nodes in cell cell 'NAND_sim{lay}'
vdd vdd 0 dc 5
vin in 0 dc 0 pulse 0 5 10n 1n 
cload out 0 250fF
.tran 0 40n
.include D:\C5_models.txt
.END

*** SPICE deck for cell 4bitupdowncounter_sim{sch} from library final_project
*** Created on Tue Dec 10, 2024 17:28:54
*** Last revised on Tue Dec 10, 2024 17:40:12
*** Written on Tue Dec 10, 2024 17:40:13 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT final_project__Dflipflop FROM CELL Dflipflop{sch}
.SUBCKT final_project__Dflipflop clk D notQ Q Res
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@546 clk net@21 gnd NMOS L=0.35U W=1.75U
Mnmos@1 D net@2 net@21 gnd NMOS L=0.35U W=1.75U
Mnmos@2 net@564 net@21 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@3 net@2 clk gnd gnd NMOS L=0.35U W=1.75U
Mnmos@4 net@820 net@564 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@11 net@222 clk net@268 gnd NMOS L=0.35U W=1.75U
Mnmos@13 Q net@241 net@268 gnd NMOS L=0.35U W=1.75U
Mnmos@15 Q notQ gnd gnd NMOS L=0.35U W=1.75U
Mnmos@16 net@222 net@564 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@22 notQ Res net@606 gnd NMOS L=0.35U W=1.75U
Mnmos@23 net@606 net@268 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@25 net@241 clk gnd gnd NMOS L=0.35U W=1.75U
Mnmos@26 net@546 Res net@820 gnd NMOS L=0.35U W=1.75U
Mpmos@0 net@21 net@2 net@546 vdd PMOS L=0.35U W=3.5U
Mpmos@1 net@21 clk D vdd PMOS L=0.35U W=3.5U
Mpmos@2 net@564 net@21 vdd vdd PMOS L=0.35U W=3.5U
Mpmos@3 net@2 clk vdd vdd PMOS L=0.35U W=3.5U
Mpmos@4 net@546 net@564 vdd vdd PMOS L=0.35U W=3.5U
Mpmos@11 net@268 net@241 net@222 vdd PMOS L=0.35U W=3.5U
Mpmos@12 net@241 clk vdd vdd PMOS L=0.35U W=3.5U
Mpmos@13 net@268 clk Q vdd PMOS L=0.35U W=3.5U
Mpmos@15 Q notQ vdd vdd PMOS L=0.35U W=3.5U
Mpmos@16 net@222 net@564 vdd vdd PMOS L=0.35U W=3.5U
Mpmos@20 net@546 Res vdd vdd PMOS L=0.35U W=3.5U
Mpmos@21 notQ Res vdd vdd PMOS L=0.35U W=3.5U
Mpmos@22 notQ net@268 vdd vdd PMOS L=0.35U W=3.5U
.ENDS final_project__Dflipflop

*** SUBCIRCUIT final_project__two_one_mux FROM CELL two_one_mux{sch}
.SUBCKT final_project__two_one_mux I0 I1 out S
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 I0 net@19 out gnd NMOS L=0.35U W=1.75U
Mnmos@1 I1 S out gnd NMOS L=0.35U W=1.75U
Mnmos@2 net@19 S gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 out S I0 vdd PMOS L=0.35U W=3.5U
Mpmos@1 out net@19 I1 vdd PMOS L=0.35U W=3.5U
Mpmos@2 net@19 S vdd vdd PMOS L=0.35U W=3.5U
.ENDS final_project__two_one_mux

*** SUBCIRCUIT final_project__4bit_up_down_counter FROM CELL 4bit_up_down_counter{sch}
.SUBCKT final_project__4bit_up_down_counter clk Q0 Q1 Q2 Q3 Res S
** GLOBAL gnd
** GLOBAL vdd
XDflipflo@0 clk net@43 net@43 Q0 Res final_project__Dflipflop
XDflipflo@1 net@9 net@52 net@52 Q1 Res final_project__Dflipflop
XDflipflo@2 net@28 net@65 net@65 Q2 Res final_project__Dflipflop
XDflipflo@3 net@12 net@75 net@75 Q3 Res final_project__Dflipflop
Xtwo_one_@0 Q0 net@43 net@9 S final_project__two_one_mux
Xtwo_one_@1 Q2 net@65 net@12 S final_project__two_one_mux
Xtwo_one_@2 Q1 net@52 net@28 S final_project__two_one_mux
.ENDS final_project__4bit_up_down_counter

.global gnd vdd

*** TOP LEVEL CELL: 4bitupdowncounter_sim{sch}
X_4bit_up_@0 clk Q0 Q1 Q2 Q3 Res S final_project__4bit_up_down_counter

* Spice Code nodes in cell cell '4bitupdowncounter_sim{sch}'
* Power Supply
vdd vdd 0 DC 3.3V
* Clock signal (50% duty cycle, period = 50ns)
vclk clk 0 PULSE(0 5 10n 1n 1n 25n 50n)
* Reset signal (Res high after first clock period)
vres res 0 PULSE(1 0 0n 5n 5n 50n 450n)
* Up-Down Select Signal (DOWN for first 200ns, then UP for remaining time)
vs s 0 PULSE(0 5 0n 1n 1n 200n 400n)
* Simulation Command
.tran 1n 450n 0 1n
* Include the D Flip-Flop and MUX Models
.include D:\C5_models.txt
.END

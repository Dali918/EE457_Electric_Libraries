*** SPICE deck for cell inverter_sim{lay} from library project_1
*** Created on Tue Oct 15, 2024 18:00:51
*** Last revised on Thu Oct 17, 2024 13:47:34
*** Written on Thu Oct 17, 2024 13:51:33 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project_1__inv_10_10 FROM CELL inv_10_10{lay}
.SUBCKT project_1__inv_10_10 gnd in out vdd
Mnmos@1 out in gnd gnd NMOS L=0.35U W=1.75U AS=4.9P AD=1.838P PS=14.35U PD=5.6U
Mpmos@1 vdd in out vdd PMOS L=0.35U W=1.75U AS=1.838P AD=4.9P PS=5.6U PD=14.35U
.ENDS project_1__inv_10_10

*** TOP LEVEL CELL: inverter_sim{lay}
Xinv_20_1@0 gnd in out vdd project_1__inv_10_10

* Spice Code nodes in cell cell 'inverter_sim{lay}'
vdd vdd 0 DC 5
vin in 0 DC 0 
.dc vin 0 5 1m
.include D:\C5_models.txt
.END

*** SPICE deck for cell inv_20_10{sch} from library tutorial_3
*** Created on Tue Oct 15, 2024 01:52:53
*** Last revised on Tue Oct 15, 2024 17:52:23
*** Written on Tue Oct 15, 2024 17:52:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inv_20_10{sch}
Mnmos@0 out in gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 out in vdd vdd PMOS L=0.35U W=3.5U

* Spice Code nodes in cell cell 'inv_20_10{sch}'
vdd vdd 0 DC 5
vin in 0 DC 0 
.dc vin 0 5 1m
.include D:\C5_models.txt
.END

*** SPICE deck for cell 8bit_ripple_bus{sch} from library project_1
*** Created on Mon Oct 21, 2024 23:29:16
*** Last revised on Mon Oct 21, 2024 23:32:15
*** Written on Mon Oct 21, 2024 23:32:20 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT project_1__full_adder FROM CELL full_adder{sch}
.SUBCKT project_1__full_adder A B Cin Cout Sout
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@17 Cin net@31 gnd NMOS L=0.35U W=1.75U
Mnmos@1 net@31 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@2 net@31 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@3 net@17 A net@30 gnd NMOS L=0.35U W=1.75U
Mnmos@4 net@30 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@5 net@108 net@17 net@125 gnd NMOS L=0.35U W=1.75U
Mnmos@6 net@125 Cin gnd gnd NMOS L=0.35U W=1.75U
Mnmos@7 net@125 B gnd gnd NMOS L=0.35U W=1.75U
Mnmos@8 net@125 A gnd gnd NMOS L=0.35U W=1.75U
Mnmos@9 net@108 A net@264 gnd NMOS L=0.35U W=1.75U
Mnmos@10 net@264 B net@263 gnd NMOS L=0.35U W=1.75U
Mnmos@11 net@263 Cin gnd gnd NMOS L=0.35U W=1.75U
Mnmos@12 Cout net@17 gnd gnd NMOS L=0.35U W=1.75U
Mnmos@13 Sout net@108 gnd gnd NMOS L=0.35U W=1.75U
Mpmos@0 net@6 Cin vdd vdd PMOS L=0.35U W=1.75U
Mpmos@1 net@83 A vdd vdd PMOS L=0.35U W=1.75U
Mpmos@2 net@6 B net@83 vdd PMOS L=0.35U W=1.75U
Mpmos@3 net@17 B net@6 vdd PMOS L=0.35U W=1.75U
Mpmos@4 net@17 A net@6 vdd PMOS L=0.35U W=1.75U
Mpmos@5 net@98 net@17 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@9 net@108 B net@98 vdd PMOS L=0.35U W=1.75U
Mpmos@10 net@108 Cin net@98 vdd PMOS L=0.35U W=1.75U
Mpmos@11 net@108 A net@98 vdd PMOS L=0.35U W=1.75U
Mpmos@12 net@205 B vdd vdd PMOS L=0.35U W=1.75U
Mpmos@13 net@207 Cin net@205 vdd PMOS L=0.35U W=1.75U
Mpmos@14 net@98 A net@207 vdd PMOS L=0.35U W=1.75U
Mpmos@15 Cout net@17 vdd vdd PMOS L=0.35U W=1.75U
Mpmos@16 Sout net@108 vdd vdd PMOS L=0.35U W=1.75U
.ENDS project_1__full_adder

.global gnd vdd

*** TOP LEVEL CELL: 8bit_ripple_bus{sch}
Xfull_add@0 full_add@0_A full_add@0_B full_add@0_Cin full_add@0_Cout full_add@0_Sout project_1__full_adder

* Spice Code nodes in cell cell '8bit_ripple_bus{sch}'
vdd vdd 0 DC 5
Va A 0 pulse 5 0 2n 1n 1n 11n 40n
Vb B 0 pulse 0 5 8n .5n .5n 8n 50n
Vc Cin 0 pulse 5 0 5n 0 0 5n 10n
.tran 20n
.include D:\C5_models.txt
.END

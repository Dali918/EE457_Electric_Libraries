*** SPICE deck for cell PMOS_IV{sch} from library tutorial_2
*** Created on Mon Oct 14, 2024 17:14:55
*** Last revised on Tue Oct 15, 2024 01:05:24
*** Written on Tue Oct 15, 2024 01:07:54 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*** WARNING: no power connection for P-transistor wells in cell 'PMOS_IV{sch}'

*** TOP LEVEL CELL: PMOS_IV{sch}
Mpmos-4@0 d g s w PMOS L=0.35U W=1.75U

* Spice Code nodes in cell cell 'PMOS_IV{sch}'
vs s 0 DC 0
vw w 0 DC 0
vg g 0 DC 0 
vd d 0 DC 0
.dc vd 0 -5 -1m vg 0 -5 -1
.include D:\C5_models.txt
.END
